

module ConnectionBox1(
	SRAM,i,o,s
);

input [0:7] SRAM;

input [0:3] i;
output [0:3] o;

input [0:3] s;


endmodule
